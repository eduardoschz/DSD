library verilog;
use verilog.vl_types.all;
entity ES201917EL_vlg_vec_tst is
end ES201917EL_vlg_vec_tst;
