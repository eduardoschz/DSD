library verilog;
use verilog.vl_types.all;
entity matrix_vlg_vec_tst is
end matrix_vlg_vec_tst;
